library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_ln2e0 is
	generic(
		word_bits	:natural:=9;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_ln2e0 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"111100011",
		"111010011",
		"111000011",
		"110110100",
		"110100110",
		"110011000",
		"110001011",
		"101111111",
		"101110011",
		"101101000",
		"101011101",
		"101010011",
		"101001001",
		"100111111",
		"100110110",
		"100101101",
		"100100101",
		"100011100",
		"100010101",
		"100001101",
		"100000110",
		"011111111",
		"011111000",
		"011110010",
		"011101100",
		"011100110",
		"011100000",
		"011011010",
		"011010101",
		"011010000",
		"011001011",
		"011000110",
		"011000001",
		"010111101",
		"010111000",
		"010110100",
		"010110000",
		"010101100",
		"010101000",
		"010100100",
		"010100001",
		"010011101",
		"010011010",
		"010010110",
		"010010011",
		"010010000",
		"010001101",
		"010001010",
		"010000111",
		"010000101",
		"010000010",
		"001111111",
		"001111101",
		"001111010",
		"001111000",
		"001110110",
		"001110011",
		"001110001",
		"001101111",
		"001101101",
		"001101011",
		"001101001",
		"001100111",
		"001100101"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)))&"000";
end architecture;