library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_reci_sqrt_1_2 is
	generic(
		word_bits	:natural:=9;
		bus_bits	:natural:=14;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_reci_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"101111100",
		"101110100",
		"101101101",
		"101100110",
		"101100000",
		"101011001",
		"101010011",
		"101001101",
		"101000110",
		"101000001",
		"100111011",
		"100110101",
		"100110000",
		"100101010",
		"100100101",
		"100100000",
		"100011011",
		"100010110",
		"100010010",
		"100001101",
		"100001000",
		"100000100",
		"100000000",
		"011111011",
		"011110111",
		"011110011",
		"011101111",
		"011101100",
		"011101000",
		"011100100",
		"011100001",
		"011011101",
		"011011010",
		"011010110",
		"011010011",
		"011010000",
		"011001101",
		"011001010",
		"011000110",
		"011000100",
		"011000001",
		"010111110",
		"010111011",
		"010111000",
		"010110110",
		"010110011",
		"010110000",
		"010101110",
		"010101011",
		"010101001",
		"010100111",
		"010100100",
		"010100010",
		"010100000",
		"010011110",
		"010011100",
		"010011001",
		"010010111",
		"010010101",
		"010010011",
		"010010001",
		"010001111",
		"010001110",
		"010001100",
		"010001010",
		"010001000",
		"010000110",
		"010000101",
		"010000011",
		"010000001",
		"010000000",
		"001111110",
		"001111101",
		"001111011",
		"001111001",
		"001111000",
		"001110111",
		"001110101",
		"001110100",
		"001110010",
		"001110001",
		"001110000",
		"001101110",
		"001101101",
		"001101100",
		"001101010",
		"001101001",
		"001101000",
		"001100111",
		"001100110",
		"001100100",
		"001100011",
		"001100010",
		"001100001",
		"001100000",
		"001011111",
		"001011110",
		"001011101",
		"001011100",
		"001011011",
		"001011010",
		"001011001",
		"001011000",
		"001010111",
		"001010110",
		"001010101",
		"001010100",
		"001010011",
		"001010010",
		"001010001",
		"001010001",
		"001010000",
		"001001111",
		"001001110",
		"001001101",
		"001001100",
		"001001100",
		"001001011",
		"001001010",
		"001001001",
		"001001001",
		"001001000",
		"001000111",
		"001000110",
		"001000110",
		"001000101",
		"001000100",
		"001000100"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)))&"000";
end architecture;