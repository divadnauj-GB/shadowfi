library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_ln2 is
	generic(
		word_bits	:natural:=16;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_ln2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"1011100010101001",
		"1011011100111011",
		"1011010111010010",
		"1011010001101111",
		"1011001100010001",
		"1011000110111000",
		"1011000001100101",
		"1010111100010110",
		"1010110111001100",
		"1010110010001000",
		"1010101101001000",
		"1010101000001100",
		"1010100011010101",
		"1010011110100011",
		"1010011001110100",
		"1010010101001011",
		"1010010000100101",
		"1010001100000011",
		"1010000111100101",
		"1010000011001011",
		"1001111110110101",
		"1001111010100011",
		"1001110110010100",
		"1001110010001001",
		"1001101110000001",
		"1001101001111101",
		"1001100101111100",
		"1001100001111111",
		"1001011110000100",
		"1001011010001101",
		"1001010110011001",
		"1001010010101000",
		"1001001110111011",
		"1001001011010000",
		"1001000111101000",
		"1001000100000011",
		"1001000000100000",
		"1000111101000001",
		"1000111001100100",
		"1000110110001001",
		"1000110010110010",
		"1000101111011101",
		"1000101100001010",
		"1000101000111010",
		"1000100101101100",
		"1000100010100001",
		"1000011111011000",
		"1000011100010001",
		"1000011001001101",
		"1000010110001010",
		"1000010011001010",
		"1000010000001100",
		"1000001101010001",
		"1000001010010111",
		"1000000111011111",
		"1000000100101001",
		"1000000001110110",
		"0111111111000100",
		"0111111100010100",
		"0111111001100110",
		"0111110110111010",
		"0111110100010000",
		"0111110001100111",
		"0111101111000000",
		"0111101100011011",
		"0111101001111000",
		"0111100111010111",
		"0111100100110111",
		"0111100010011000",
		"0111011111111100",
		"0111011101100000",
		"0111011011000111",
		"0111011000101111",
		"0111010110011000",
		"0111010100000011",
		"0111010001110000",
		"0111001111011110",
		"0111001101001101",
		"0111001010111110",
		"0111001000110000",
		"0111000110100011",
		"0111000100011000",
		"0111000010001110",
		"0111000000000110",
		"0110111101111110",
		"0110111011111000",
		"0110111001110100",
		"0110110111110000",
		"0110110101101110",
		"0110110011101101",
		"0110110001101101",
		"0110101111101110",
		"0110101101110000",
		"0110101011110100",
		"0110101001111001",
		"0110100111111110",
		"0110100110000101",
		"0110100100001101",
		"0110100010010110",
		"0110100000100000",
		"0110011110101011",
		"0110011100110111",
		"0110011011000101",
		"0110011001010011",
		"0110010111100010",
		"0110010101110010",
		"0110010100000011",
		"0110010010010101",
		"0110010000101000",
		"0110001110111011",
		"0110001101010000",
		"0110001011100110",
		"0110001001111100",
		"0110001000010100",
		"0110000110101100",
		"0110000101000101",
		"0110000011011111",
		"0110000001111010",
		"0110000000010101",
		"0101111110110010",
		"0101111101001111",
		"0101111011101101",
		"0101111010001100",
		"0101111000101011",
		"0101110111001100",
		"0101110101101101",
		"0101110100001111",
		"0101110010110001"
	);
begin
	data <= "0"&rom(to_integer(unsigned(addr)))&"000";
end architecture;