module dummy;

endmodule;