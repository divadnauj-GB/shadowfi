library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_sqrt_2_4 is
	generic(
		word_bits	:natural:=25;
		bus_bits	:natural:=29;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"0110101000001001111001101",
		"0110110011011011001010111",
		"0110111110100110111010100",
		"0111001001101101010000011",
		"0111010100101110010100010",
		"0111011111101010001101011",
		"0111101010100001000011010",
		"0111110101010010111100100",
		"1000000000000000000000000",
		"1000001010101000010100000",
		"1000010101001011111110110",
		"1000011111101011000110011",
		"1000101010000101110000100",
		"1000110100011100000011000",
		"1000111110101110000011000",
		"1001001000111011110101111",
		"1001010011000101100000111",
		"1001011101001011001000110",
		"1001100111001100110010011",
		"1001110001001010100010010",
		"1001111011000100011101001",
		"1010000100111010100111001",
		"1010001110101101000100101",
		"1010011000011011111001101",
		"1010100010000111001010010",
		"1010101011101110111010011",
		"1010110101010011001101101",
		"1010111110110100000111110",
		"1011001000010001101100011",
		"1011010001101011111111000",
		"1011011011000011000010111",
		"1011100100010110111011010",
		"1011101101100111101011101",
		"1011110110110101010110110",
		"1100000000000000000000000",
		"1100001001000111101010000",
		"1100010010001100011000000",
		"1100011011001110001100100",
		"1100100100001101001010011",
		"1100101101001001010100011",
		"1100110110000010101101000",
		"1100111110111001010110111",
		"1101000111101101010100100",
		"1101010000011110101000001",
		"1101011001001101010100011",
		"1101100001111001011011100",
		"1101101010100010111111110",
		"1101110011001010000011010",
		"1101111011101110101000010",
		"1110000100010000110000111",
		"1110001100110000011111001",
		"1110010101001101110101001",
		"1110011101101000110100111",
		"1110100110000001100000001",
		"1110101110010111111001000",
		"1110110110101100000001010",
		"1110111110111101111010110",
		"1111000111001101100111001",
		"1111001111011011001000010",
		"1111010111100110011111111",
		"1111011111101111101111101",
		"1111100111110110111001001",
		"1111101111111011111101111",
		"1111110111111110111111110"
	);
begin
	data <= "01"&rom(to_integer(unsigned(addr)))&"00";
end architecture;