library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_exp is
	generic(
		word_bits	:natural:=16;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_exp is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"0101100010111000",
		"0101100110110000",
		"0101101010101010",
		"0101101110100110",
		"0101110010100110",
		"0101110110101000",
		"0101111010101101",
		"0101111110110101",
		"0110000011000000",
		"0110000111001110",
		"0110001011011110",
		"0110001111110010",
		"0110010100001001",
		"0110011000100010",
		"0110011100111111",
		"0110100001011111",
		"0110100110000010",
		"0110101010101000",
		"0110101111010001",
		"0110110011111110",
		"0110111000101110",
		"0110111101100001",
		"0111000010010111",
		"0111000111010001",
		"0111001100001110",
		"0111010001001111",
		"0111010110010011",
		"0111011011011011",
		"0111100000100110",
		"0111100101110101",
		"0111101011001000",
		"0111110000011110",
		"0111110101111000",
		"0111111011010110",
		"1000000000111000",
		"1000000110011101",
		"1000001100000110",
		"1000010001110100",
		"1000010111100101",
		"1000011101011010",
		"1000100011010011",
		"1000101001010001",
		"1000101111010010",
		"1000110101011000",
		"1000111011100010",
		"1001000001110001",
		"1001001000000011",
		"1001001110011010",
		"1001010100110110",
		"1001011011010110",
		"1001100001111010",
		"1001101000100011",
		"1001101111010001",
		"1001110110000011",
		"1001111100111010",
		"1010000011110110",
		"1010001010110111",
		"1010010001111101",
		"1010011001000111",
		"1010100000010111",
		"1010100111101011",
		"1010101111000101",
		"1010110110100100",
		"1010111110001000"
	);
begin
	data <= "0"&rom(to_integer(unsigned(addr)))&"000";
end architecture;