library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_ln2e0 is
	generic(
		word_bits	:natural:=25;
		bus_bits	:natural:=29;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_ln2e0 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"1110001010101000111010110",
		"1101110011110010110011110",
		"1101011101011010011011010",
		"1101000111011110110001000",
		"1100110001111110110111100",
		"1100011100111001110100100",
		"1100001000001110110000010",
		"1011110011111100110101100",
		"1011100000000011010001100",
		"1011001100100001010011110",
		"1010111001010110001101101",
		"1010100110100001010010111",
		"1010010100000001111000111",
		"1010000001110111010110111",
		"1001110000000001000101111",
		"1001011110011110100000010",
		"1001001101001111000010001",
		"1000111100010010001001000",
		"1000101011100111010011110",
		"1000011011001110000010011",
		"1000001011000101110110011",
		"0111111011001110010010011",
		"0111101011100110111001110",
		"0111011100001111010001100",
		"0111001101000110111111001",
		"0110111110001101101001100",
		"0110101111100010111000000",
		"0110100001000110010011010",
		"0110010010110111100100011",
		"0110000100110110010101110",
		"0101110111000010010001111",
		"0101101001011011000100101",
		"0101011100000000011010001",
		"0101001110110001111111010",
		"0101000001101111100001101",
		"0100110100111000101111011",
		"0100101000001101010111010",
		"0100011011101101001000110",
		"0100001111010111110011011",
		"0100000011001101000111110",
		"0011110111001100110110101",
		"0011101011010110110001010",
		"0011011111101010101001100",
		"0011010100001000010001101",
		"0011001000101111011100000",
		"0010111101011111111011111",
		"0010110010011001100100100",
		"0010100111011100001001110",
		"0010011100100111011111111",
		"0010010001111011011011000",
		"0010000111010111110000011",
		"0001111100111100010100110",
		"0001110010101000111101110",
		"0001101000011101100001000",
		"0001011110011001110100101",
		"0001010100011101101111000",
		"0001001010101001000110011",
		"0001000000111011110001111",
		"0000110111010101101000011",
		"0000101101110110100001010",
		"0000100100011110010100000",
		"0000011011001100111000011",
		"0000010010000010000110010",
		"0000001000111101110110000"
	);
begin
	data <= "010"&rom(to_integer(unsigned(addr)))&"0";
end architecture;