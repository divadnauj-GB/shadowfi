library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_ln2 is
	generic(
		word_bits	:natural:=26;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_ln2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"00000000000000000000000000",
		"00000010110111111100101000",
		"00000101101110011110010110",
		"00001000100011100110100100",
		"00001011010111010110100111",
		"00001110001001101111110101",
		"00010000111010110011100010",
		"00010011101010100010111111",
		"00010110011000111111011100",
		"00011001000110001010000110",
		"00011011110010000100001001",
		"00011110011100101110110000",
		"00100001000110001011000100",
		"00100011101110011010001101",
		"00100110010101011101001111",
		"00101000111011010101010000",
		"00101011100000000011010010",
		"00101110000011101000010110",
		"00110000100110000101011110",
		"00110011000111011011101000",
		"00110101100111101011110001",
		"00111000000110110110110110",
		"00111010100100111101110010",
		"00111101000010000001011111",
		"00111111011110000010110110",
		"01000001111001000010101110",
		"01000100010011000001111101",
		"01000110101100000001011011",
		"01001001000100000001111010",
		"01001011011011000100010000",
		"01001101110001001001001101",
		"01010000000110010001100011",
		"01010010011010011110000100",
		"01010100101101101111100000",
		"01010111000000000110100011",
		"01011001010001100011111110",
		"01011011100010001000011101",
		"01011101110001110100101011",
		"01100000000000101001010110",
		"01100010001110100111000111",
		"01100100011011101110101000",
		"01100110101000000000100011",
		"01101000110011011101100000",
		"01101010111110000110000111",
		"01101101000111111010111111",
		"01101111010000111100101110",
		"01110001011001001011111011",
		"01110011100000101001001001",
		"01110101100111010100111110",
		"01110111101101001111111101",
		"01111001110010011010101010",
		"01111011110110110101100111",
		"01111101111010100001010110",
		"01111111111101011110011001",
		"10000001111111101101010001",
		"10000100000001001110011110",
		"10000110000010000010100000",
		"10001000000010001001110110",
		"10001010000001100100111111",
		"10001100000000010100011010",
		"10001101111110011000100011",
		"10001111111011110001111010",
		"10010001111000100000111010",
		"10010011110100100110000000",
		"10010101110000000001101001",
		"10010111101010110100001110",
		"10011001100100111110001101",
		"10011011011110011111111111",
		"10011101010111011001111111",
		"10011111001111101100100111",
		"10100001000111011000001111",
		"10100010111110011101010011",
		"10100100110100111100001001",
		"10100110101010110101001011",
		"10101000100000001000110001",
		"10101010010100110111010001",
		"10101100001001000001000100",
		"10101101111100100110100001",
		"10101111101111100111111110",
		"10110001100010000101110010",
		"10110011010100000000010001",
		"10110101000101010111110011",
		"10110110110110001100101101",
		"10111000100110011111010011",
		"10111010010110001111111010",
		"10111100000101011110111000",
		"10111101110100001100011111",
		"10111111100010011001000100",
		"11000001010000000100111010",
		"11000010111101010000010110",
		"11000100101001111011101001",
		"11000110010110000111000111",
		"11001000000001110011000010",
		"11001001101100111111101101",
		"11001011010111101101011010",
		"11001101000001111100011010",
		"11001110101011101100111111",
		"11010000010100111111011011",
		"11010001111101110011111110",
		"11010011100110001010111010",
		"11010101001110000100011110",
		"11010110110101100000111100",
		"11011000011100100000100100",
		"11011010000011000011100110",
		"11011011101001001010010010",
		"11011101001110110100110110",
		"11011110110100000011100011",
		"11100000011000110110101000",
		"11100001111101001110010100",
		"11100011100001001010110101",
		"11100101000100101100011011",
		"11100110100111110011010100",
		"11101000001010011111101101",
		"11101001101100110001110110",
		"11101011001110101001111100",
		"11101100110000001000001100",
		"11101110010001001100110101",
		"11101111110001111000000100",
		"11110001010010001010000101",
		"11110010110010000011000111",
		"11110100010001100011010110",
		"11110101110000101010111111",
		"11110111001111011010001110",
		"11111000101101110001010000",
		"11111010001011110000010001",
		"11111011101001010111011110",
		"11111101000110100111000010",
		"11111110100011011111001001"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)))&"0";
end architecture;