library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_reci_sqrt_2_4 is
	generic(
		word_bits	:natural:=9;
		bus_bits	:natural:=14;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_reci_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"100001100",
		"100000111",
		"100000010",
		"011111101",
		"011111001",
		"011110100",
		"011101111",
		"011101011",
		"011100111",
		"011100011",
		"011011110",
		"011011010",
		"011010111",
		"011010011",
		"011001111",
		"011001100",
		"011001000",
		"011000101",
		"011000001",
		"010111110",
		"010111011",
		"010111000",
		"010110101",
		"010110010",
		"010101111",
		"010101100",
		"010101001",
		"010100110",
		"010100100",
		"010100001",
		"010011111",
		"010011100",
		"010011010",
		"010010111",
		"010010101",
		"010010011",
		"010010001",
		"010001110",
		"010001100",
		"010001010",
		"010001000",
		"010000110",
		"010000100",
		"010000010",
		"010000000",
		"001111110",
		"001111101",
		"001111011",
		"001111001",
		"001110111",
		"001110110",
		"001110100",
		"001110010",
		"001110001",
		"001101111",
		"001101110",
		"001101100",
		"001101011",
		"001101001",
		"001101000",
		"001100111",
		"001100101",
		"001100100",
		"001100011",
		"001100001",
		"001100000",
		"001011111",
		"001011110",
		"001011100",
		"001011011",
		"001011010",
		"001011001",
		"001011000",
		"001010111",
		"001010110",
		"001010101",
		"001010100",
		"001010011",
		"001010010",
		"001010001",
		"001010000",
		"001001111",
		"001001110",
		"001001101",
		"001001100",
		"001001011",
		"001001010",
		"001001001",
		"001001000",
		"001001000",
		"001000111",
		"001000110",
		"001000101",
		"001000100",
		"001000100",
		"001000011",
		"001000010",
		"001000001",
		"001000001",
		"001000000",
		"000111111",
		"000111111",
		"000111110",
		"000111101",
		"000111101",
		"000111100",
		"000111011",
		"000111011",
		"000111010",
		"000111001",
		"000111001",
		"000111000",
		"000111000",
		"000110111",
		"000110110",
		"000110110",
		"000110101",
		"000110101",
		"000110100",
		"000110100",
		"000110011",
		"000110011",
		"000110010",
		"000110010",
		"000110001",
		"000110001",
		"000110000",
		"000110000"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)))&"000";
end architecture;