library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_sqrt_1_2 is
	generic(
		word_bits	:natural:=13;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"1111111111111",
		"1111110000001",
		"1111100000101",
		"1111010001100",
		"1111000010110",
		"1110110100010",
		"1110100110001",
		"1110011000011",
		"1110001010110",
		"1101111101100",
		"1101110000100",
		"1101100011110",
		"1101010111010",
		"1101001011000",
		"1100111111000",
		"1100110011010",
		"1100100111110",
		"1100011100011",
		"1100010001010",
		"1100000110010",
		"1011111011100",
		"1011110001000",
		"1011100110101",
		"1011011100100",
		"1011010010100",
		"1011001000101",
		"1010111111000",
		"1010110101011",
		"1010101100001",
		"1010100010111",
		"1010011001110",
		"1010010000111",
		"1010001000001",
		"1001111111100",
		"1001110111000",
		"1001101110101",
		"1001100110011",
		"1001011110010",
		"1001010110001",
		"1001001110010",
		"1001000110100",
		"1000111110111",
		"1000110111010",
		"1000101111111",
		"1000101000100",
		"1000100001010",
		"1000011010001",
		"1000010011000",
		"1000001100001",
		"1000000101010",
		"0111111110011",
		"0111110111110",
		"0111110001001",
		"0111101010101",
		"0111100100010",
		"0111011101111",
		"0111010111101",
		"0111010001011",
		"0111001011010",
		"0111000101010",
		"0110111111010",
		"0110111001011",
		"0110110011100",
		"0110101101110"
	);
begin
	data <= "0001"&rom(to_integer(unsigned(addr)))&"000";
end architecture;