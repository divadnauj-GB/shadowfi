library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_reci is
	generic(
		word_bits	:natural:=16;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_reci is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"1111111111111101",
		"1111110000001001",
		"1111100000101100",
		"1111010001100110",
		"1111000010110110",
		"1110110100011011",
		"1110100110010100",
		"1110011000100010",
		"1110001011000010",
		"1101111101110110",
		"1101110000111100",
		"1101100100010100",
		"1101010111111101",
		"1101001011110110",
		"1101000000000000",
		"1100110100011010",
		"1100101001000100",
		"1100011101111100",
		"1100010011000011",
		"1100001000011000",
		"1011111101111011",
		"1011110011101011",
		"1011101001101000",
		"1011011111110010",
		"1011010110001001",
		"1011001100101011",
		"1011000011011001",
		"1010111010010011",
		"1010110001011000",
		"1010101000101000",
		"1010100000000010",
		"1010010111100111",
		"1010001111010110",
		"1010000111001110",
		"1001111111010000",
		"1001110111011100",
		"1001101111110001",
		"1001101000001110",
		"1001100000110101",
		"1001011001100011",
		"1001010010011010",
		"1001001011011001",
		"1001000100100000",
		"1000111101101111",
		"1000110111000101",
		"1000110000100011",
		"1000101010001000",
		"1000100011110100",
		"1000011101100111",
		"1000010111100000",
		"1000010001100000",
		"1000001011100110",
		"1000000101110011",
		"1000000000000110",
		"0111111010011111",
		"0111110100111101",
		"0111101111100010",
		"0111101010001100",
		"0111100100111100",
		"0111011111110001",
		"0111011010101011",
		"0111010101101010",
		"0111010000101111",
		"0111001011111000",
		"0111000111000110",
		"0111000010011001",
		"0110111101110001",
		"0110111001001101",
		"0110110100101101",
		"0110110000010010",
		"0110101011111100",
		"0110100111101001",
		"0110100011011011",
		"0110011111010000",
		"0110011011001010",
		"0110010111000111",
		"0110010011001000",
		"0110001111001101",
		"0110001011010110",
		"0110000111100010",
		"0110000011110010",
		"0110000000000101",
		"0101111100011011",
		"0101111000110101",
		"0101110101010010",
		"0101110001110010",
		"0101101110010101",
		"0101101010111100",
		"0101100111100101",
		"0101100100010010",
		"0101100001000001",
		"0101011101110011",
		"0101011010101000",
		"0101010111100000",
		"0101010100011010",
		"0101010001010111",
		"0101001110010111",
		"0101001011011001",
		"0101001000011110",
		"0101000101100101",
		"0101000010101111",
		"0100111111111011",
		"0100111101001001",
		"0100111010011010",
		"0100110111101100",
		"0100110101000010",
		"0100110010011001",
		"0100101111110010",
		"0100101101001110",
		"0100101010101100",
		"0100101000001011",
		"0100100101101101",
		"0100100011010001",
		"0100100000110110",
		"0100011110011110",
		"0100011100000111",
		"0100011001110010",
		"0100010111100000",
		"0100010101001110",
		"0100010010111111",
		"0100010000110001",
		"0100001110100101",
		"0100001100011011",
		"0100001010010011",
		"0100001000001100",
		"0100000110000110",
		"0100000100000010",
		"0100000010000000"
	);
begin
	data <= "10"&rom(to_integer(unsigned(addr)))&"00";
end architecture;