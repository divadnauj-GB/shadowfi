library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_sqrt_1_2 is
	generic(
		word_bits	:natural:=8;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"11111101",
		"11110111",
		"11110001",
		"11101100",
		"11100111",
		"11100010",
		"11011101",
		"11011000",
		"11010100",
		"11010000",
		"11001011",
		"11000111",
		"11000011",
		"11000000",
		"10111100",
		"10111000",
		"10110101",
		"10110010",
		"10101110",
		"10101011",
		"10101000",
		"10100101",
		"10100010",
		"10100000",
		"10011101",
		"10011010",
		"10011000",
		"10010101",
		"10010011",
		"10010000",
		"10001110",
		"10001100",
		"10001010",
		"10001000",
		"10000110",
		"10000100",
		"10000010",
		"10000000",
		"01111110",
		"01111100",
		"01111010",
		"01111000",
		"01110111",
		"01110101",
		"01110011",
		"01110010",
		"01110000",
		"01101111",
		"01101101",
		"01101100",
		"01101010",
		"01101001",
		"01101000",
		"01100110",
		"01100101",
		"01100100",
		"01100011",
		"01100001",
		"01100000",
		"01011111",
		"01011110",
		"01011101",
		"01011100",
		"01011011"
	);
begin
	data <= "1000"&rom(to_integer(unsigned(addr)))&"00";
end architecture;